`include "opcodes.v"
`include "alu_opcodes.v"

module ALU(input [4:0] alu_op,
           input [31:0] alu_in_1,
           input [31:0] alu_in_2,      
           output [31:0] alu_result,        
           output alu_bcond);  
endmodule
