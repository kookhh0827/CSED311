`include "opcodes.v"
`include "alu_opcodes.v"

module ImmediateGenerator(input [31:0] instr,   
                          output [31:0] imm_gen_out);  
endmodule
