module ALUControlUnit(input [6:0] opcode,
                      input [2:0] funct3,
                      input [6:0] funct7,      
                      output [8:0] alu_op);  
endmodule
