module AddressSelector(input [6:0] opcode,
                       input cs_plus_1,
                       input [1:0] AddrCtl,
                       input alu_bcond,
                       input ns_IF1,
                       input is_ecall,
                       output reg [4:0] next_state);
    
endmodule

